netcdf test_1d_arrays {
// Global attributes

group: testGroup {

dimensions:
    arraysize = 3;

variables:
    byte simpleByte(arraysize);
    short simpleShort(arraysize);
    int simpleInt(arraysize);
    float simpleFloat(arraysize);
    double simpleDouble(arraysize);

data:
   
   simpleByte = 1,2,3;
   simpleShort = 1,2,3;
   simpleInt = 1,2,3;
   simpleFloat = 4.5,5.5,6.6;
   simpleDouble = 4.5,5.5,6.6;
}
}
