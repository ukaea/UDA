netcdf test_string {
// Global attributes

group: testGroup {

variables:
    string simpleString;

data:
   
   simpleString = "Hello";
}
}
