netcdf test_compound_scalars {
// Global attributes

group: testGroup {

types:
  compound testCompoundByte {
    byte simpleByte;
  }

  compound testCompoundShort {
    int simpleShort;
  }

  compound testCompoundInt {
    int simpleInt;
  }

  compound testCompoundFloat {
    float simpleFloat;
  }

  compound testCompoundDouble {
    double simpleDouble;
  }

dimensions:
  arraySize = 2;

variables:
  testCompoundByte simpleByte(arraySize);
  testCompoundByte simpleShort(arraySize);
  testCompoundInt simpleInt(arraySize);
  testCompoundFloat simpleFloat(arraySize);
  testCompoundDouble simpleDouble(arraySize);

data:
   
   simpleByte = {1},{2};
   simpleShort = {1},{2};
   simpleInt = {1},{2};
   simpleFloat = {4.5},{4.4};
   simpleDouble = {4.5},{4.4};
}
}
