netcdf test_string_arrays {
// Global attributes

group: testGroup {

dimensions:
    arraySize = 3;

variables:
    string simpleString(arraySize);

data:
   
   simpleString = "Hello", "Hi", "Good Day";
}
}
