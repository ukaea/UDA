netcdf test_compound_nested_1d_arrays {
// Global attributes

group: testGroup {

types:

  compound testCompoundFloatScalar {
    float simpleFloat;        
  }

  compound testCompoundFloat {
    float simpleFloat(3);        
  }

  compound testCompoundFloatLonger {
    float simpleFloat(10);        
  }

  compound testCompound {
    string name;
    float something;
    testCompoundFloatScalar scalar;
    testCompoundFloat shortarray;
    testCompoundFloatLonger longarray;
  }

dimensions:
 singleDim = 1;

variables:
  testCompound simpleFloatVar(singleDim);

data:
   simpleFloatVar = {"test", 223.9, {1.0}, {{4.5,5.5,6.6}}, {{1,2,3,4,5,6,7,8,9,10}} };
}
}
