netcdf test_2d_arrays {
// Global attributes

group: testGroup {

dimensions:
    arraysize1 = 3;
    arraysize2 = 2;

variables:
    byte simpleByte(arraysize1, arraysize2);
    short simpleShort(arraysize1, arraysize2);
    int simpleInt(arraysize1, arraysize2);
    float simpleFloat(arraysize1, arraysize2);
    double simpleDouble(arraysize1, arraysize2);

data:
   
   simpleByte = 1,2,3, 
                1,2,3;
   simpleShort = 1,2,3, 
                 1,2,3;   
   simpleInt =  1,2,3, 
                1,2,3;
   simpleFloat = 4.5,5.5,6.6, 
                 4.5,5.5,6.6;
   simpleDouble = 4.5,5.5,6.6, 
                  4.5,5.5,6.6;
}
}
